// Code your testbench here
// or browse Examples

//`include "z_comp_tb.sv"
`include "cordic_comp_tb.sv"

// `include "counter_mod_tb.sv"

//`include "mux_input_controller_tb.sv"
// Code your design here

//`include "z_comp.sv"
`include "cordic_comp.sv"

`include "di_ei_LUT.sv"

`include "di_control_comp.sv"

`include "dff.sv"

`include "reg_2to1_mux.sv"

`include "addorsub_2to1_mux.sv"

`include "shifter.sv"

`include "counter_mod.sv"

`include "mux_input_controller.sv"
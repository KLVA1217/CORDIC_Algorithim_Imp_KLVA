// Code your design here
module di_ei_LUT
   (input  [5:0] count,
    output reg [63:0] di_ei_result);
  
  // reg [63:0] di_ei_result;
  
  always @ (count) begin
    case(count) // arctan(2^i) or tan(arctan(2^i)) in radians converted to binary
		6'b00 : di_ei_result <= 64'b0110010010000111111011010101000100010000101101000110000000000000;// arctan(2^-0)
		6'b01 : di_ei_result <= 64'b0011101101011000110011100000101011000011011101101001111000000000;// arctan(2^-1)
		6'b10 : di_ei_result <= 64'b0001111101011011011101011111100100101100100000001101110100000000;// arctan(2^-2)
		6'b11 : di_ei_result <= 64'b0000111111101010110111010100110101010110000101111011011100000000;// arctan(2^-3)
		6'b100 : di_ei_result <= 64'b0000011111111101010101101110110111001011001111110111101010000000;// arctan(2^-4)
		6'b101 : di_ei_result <= 64'b0000001111111111101010101011011101110101001011101100010010100000;// arctan(2^-5)
		6'b110 : di_ei_result <= 64'b0000000111111111111101010101010110111011101101110010100110110000;// arctan(2^-6)
		6'b111 : di_ei_result <= 64'b0000000011111111111111101010101010101101110111011101010010111000;// arctan(2^-7)
		6'b1000 : di_ei_result <= 64'b0000000001111111111111111101010101010101011011101110111011011100;// arctan(2^-8)
		6'b1001 : di_ei_result <= 64'b0000000000111111111111111111101010101010101010110111011101111000;// arctan(2^-9)
		6'b1010 : di_ei_result <= 64'b0000000000011111111111111111111101010101010101010101101110111100;// arctan(2^-10)
		6'b1011 : di_ei_result <= 64'b0000000000001111111111111111111111101010101010101010101011011110;// arctan(2^-11)
		6'b1100 : di_ei_result <= 64'b0000000000000111111111111111111111111101010101010101010101010111;// arctan(2^-12)
		6'b1101 : di_ei_result <= 64'b0000000000000011111111111111111111111111101010101010101010101010;// arctan(2^-13)
		6'b1110 : di_ei_result <= 64'b0000000000000001111111111111111111111111111101010101010101010101;// arctan(2^-14)
		6'b1111 : di_ei_result <= 64'b0000000000000000111111111111111111111111111111101010101010101010;// arctan(2^-15)
		6'b10000 : di_ei_result <= 64'b0000000000000000011111111111111111111111111111111101010101010101;// arctan(2^-16)
		6'b10001 : di_ei_result <= 64'b0000000000000000001111111111111111111111111111111111101010101010;// arctan(2^-17)
		6'b10010 : di_ei_result <= 64'b0000000000000000000111111111111111111111111111111111111101010101;// arctan(2^-18)
		6'b10011 : di_ei_result <= 64'b0000000000000000000011111111111111111111111111111111111111101010;// arctan(2^-19)
		6'b10100 : di_ei_result <= 64'b0000000000000000000001111111111111111111111111111111111111111101;// arctan(2^-20)
		6'b10101 : di_ei_result <= 64'b0000000000000000000000111111111111111111111111111111111111111111;// arctan(2^-21)
		6'b10110 : di_ei_result <= 64'b0000000000000000000000011111111111111111111111111111111111111111;// arctan(2^-22)
		6'b10111 : di_ei_result <= 64'b0000000000000000000000001111111111111111111111111111111111111111;// arctan(2^-23)
		6'b11000 : di_ei_result <= 64'b0000000000000000000000000111111111111111111111111111111111111111;// arctan(2^-24)
		6'b11001 : di_ei_result <= 64'b0000000000000000000000000011111111111111111111111111111111111111;// arctan(2^-25)
		6'b11010 : di_ei_result <= 64'b0000000000000000000000000001111111111111111111111111111111111111;// arctan(2^-26)
		6'b11011 : di_ei_result <= 64'b0000000000000000000000000001000000000000000000000000000000000000;// arctan(2^-27)
		6'b11100 : di_ei_result <= 64'b0000000000000000000000000000100000000000000000000000000000000000;// arctan(2^-28)
		6'b11101 : di_ei_result <= 64'b0000000000000000000000000000010000000000000000000000000000000000;// arctan(2^-29)
		6'b11110 : di_ei_result <= 64'b0000000000000000000000000000001000000000000000000000000000000000;// arctan(2^-30)
		6'b11111 : di_ei_result <= 64'b0000000000000000000000000000000100000000000000000000000000000000;// arctan(2^-31)
		6'b100000 : di_ei_result <= 64'b0000000000000000000000000000000010000000000000000000000000000000;// arctan(2^-32)
		6'b100001 : di_ei_result <= 64'b0000000000000000000000000000000001000000000000000000000000000000;// arctan(2^-33)
		6'b100010 : di_ei_result <= 64'b0000000000000000000000000000000000100000000000000000000000000000;// arctan(2^-34)
		6'b100011 : di_ei_result <= 64'b0000000000000000000000000000000000010000000000000000000000000000;// arctan(2^-35)
		6'b100100 : di_ei_result <= 64'b0000000000000000000000000000000000001000000000000000000000000000;// arctan(2^-36)
		6'b100101 : di_ei_result <= 64'b0000000000000000000000000000000000000100000000000000000000000000;// arctan(2^-37)
		6'b100110 : di_ei_result <= 64'b0000000000000000000000000000000000000010000000000000000000000000;// arctan(2^-38)
		6'b100111 : di_ei_result <= 64'b0000000000000000000000000000000000000001000000000000000000000000;// arctan(2^-39)
		6'b101000 : di_ei_result <= 64'b0000000000000000000000000000000000000000100000000000000000000000;// arctan(2^-40)
		6'b101001 : di_ei_result <= 64'b0000000000000000000000000000000000000000010000000000000000000000;// arctan(2^-41)
		6'b101010 : di_ei_result <= 64'b0000000000000000000000000000000000000000001000000000000000000000;// arctan(2^-42)
		6'b101011 : di_ei_result <= 64'b0000000000000000000000000000000000000000000100000000000000000000;// arctan(2^-43)
		6'b101100 : di_ei_result <= 64'b0000000000000000000000000000000000000000000010000000000000000000;// arctan(2^-44)
		6'b101101 : di_ei_result <= 64'b0000000000000000000000000000000000000000000001000000000000000000;// arctan(2^-45)
		6'b101110 : di_ei_result <= 64'b0000000000000000000000000000000000000000000000100000000000000000;// arctan(2^-46)
		6'b101111 : di_ei_result <= 64'b0000000000000000000000000000000000000000000000010000000000000000;// arctan(2^-47)
		6'b110000 : di_ei_result <= 64'b0000000000000000000000000000000000000000000000001000000000000000;// arctan(2^-48)
		6'b110001 : di_ei_result <= 64'b0000000000000000000000000000000000000000000000000100000000000000;// arctan(2^-49)
		6'b110010 : di_ei_result <= 64'b0000000000000000000000000000000000000000000000000010000000000000;// arctan(2^-50)
		6'b110011 : di_ei_result <= 64'b0000000000000000000000000000000000000000000000000001000000000000;// arctan(2^-51)
		6'b110100 : di_ei_result <= 64'b0000000000000000000000000000000000000000000000000000100000000000;// arctan(2^-52)
		6'b110101 : di_ei_result <= 64'b0000000000000000000000000000000000000000000000000000010000000000;// arctan(2^-53)
		6'b110110 : di_ei_result <= 64'b0000000000000000000000000000000000000000000000000000001000000000;// arctan(2^-54)
		6'b110111 : di_ei_result <= 64'b0000000000000000000000000000000000000000000000000000000100000000;// arctan(2^-55)
		6'b111000 : di_ei_result <= 64'b0000000000000000000000000000000000000000000000000000000010000000;// arctan(2^-56)
		6'b111001 : di_ei_result <= 64'b0000000000000000000000000000000000000000000000000000000001000000;// arctan(2^-57)
		6'b111010 : di_ei_result <= 64'b0000000000000000000000000000000000000000000000000000000000100000;// arctan(2^-58)
		6'b111011 : di_ei_result <= 64'b0000000000000000000000000000000000000000000000000000000000010000;// arctan(2^-59)
		6'b111100 : di_ei_result <= 64'b0000000000000000000000000000000000000000000000000000000000001000;// arctan(2^-60)
		6'b111101 : di_ei_result <= 64'b0000000000000000000000000000000000000000000000000000000000000100;// arctan(2^-61)
		6'b111110 : di_ei_result <= 64'b0000000000000000000000000000000000000000000000000000000000000010;// arctan(2^-62)
		6'b111111 : di_ei_result <= 64'b0000000000000000000000000000000000000000000000000000000000000001;// arctan(2^-63)
      default: di_ei_result <= 0;
    endcase
    
    //di_ei_output = di_ei_result[63 : (63 - (BIT_WIDTH - 1))];
    
  end
endmodule
// Code your testbench here
// or browse Examples

// `include "dff_tb.sv"

// `include "di_control_comp_tb.sv"

// `include "reg_2to1_mux_tb.sv"

// `include "addorsub_2to1_mux_tb.sv"

// `include "di_ei_LUT_tb.sv"

// `include "shifter_tb.sv"

// `include "counter_mod_tb.sv"

`include "cordic_comp_tb.sv"